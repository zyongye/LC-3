`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/22/2019 06:22:00 PM
// Design Name: 
// Module Name: CtrlStore
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module CtrlStore(
    input [5:0] uPC,
    output [48:0] uInstruction
    );

    reg [48:0] uInstructionStore[63:0];

    initial begin
        uInstructionStore[0] = 49'b0010010010000000000000000000000000000000000000000;
        uInstructionStore[1] = 49'b0000010010000011000000010000000000100000000000000;
        uInstructionStore[2] = 49'b0000011001100000000000001000000000001000100000000;
        uInstructionStore[3] = 49'b0000010111100000000000001000000000001000100000000;
        uInstructionStore[4] = 49'b0000010100000000000000000000000000000000000000000; 
        uInstructionStore[5] = 49'b0000010010000011000000010000000000100000000001000;
        uInstructionStore[6] = 49'b0000011001100000000000001000000000110100100000000;
        uInstructionStore[7] = 49'b0000010111100000000000001000000000110100100000000;
        uInstructionStore[9] = 49'b0000010010000011000000010000000000100000000010000;
        uInstructionStore[10] = 49'b0000011000100000000000001000000000001000100000000;
        uInstructionStore[11] = 49'b0000011101100000000000001000000000001000100000000;
        uInstructionStore[12] = 49'b0000010010000000100000000000010000110000000000000;
        uInstructionStore[14] = 49'b0000010010000011000000001000000000001000000000000;
        uInstructionStore[15] = 49'b0000011100100000000000001000000000000000000000000;
        uInstructionStore[16] = 49'b0001010000000000000000000000000000000000000000110;
        uInstructionStore[18] = 49'b0101100001100000100001000000000000000000000000000;
        uInstructionStore[20] = 49'b0000010010000010100001000000010010110000000000000;
        uInstructionStore[21] = 49'b0000010010000010100001000000010010001100000000000;
        uInstructionStore[22] = 49'b0000010010000000100000000000010000001000000000000;
        uInstructionStore[23] = 49'b0000010000010000000000010000000000000000000011000;
        uInstructionStore[24] = 49'b0001011000010000000000000000000000000000000000100;
        uInstructionStore[25] = 49'b0001011001010000000000000000000000000000000000100;
        uInstructionStore[26] = 49'b0000011001100000000000100000000000000000000000000;
        uInstructionStore[27] = 49'b0000010010000011000000100000000000000000000000000;
        uInstructionStore[28] = 49'b0001011100010010000001000000000010000000000000010;
        uInstructionStore[29] = 49'b0001011101010000000000000000000000000000000000100;
        uInstructionStore[30] = 49'b0000010010000000100000100000011000000000000000000;
        uInstructionStore[31] = 49'b0000010111100000000000100000000000000000000000000;
        uInstructionStore[32] = 49'b1000xxxxxx000100000000000000000000000000000000000;
        uInstructionStore[33] = 49'b0001100001010000000000000000000000000000000000100;
        uInstructionStore[35] = 49'b0000100000001000000000100000000000000000000000000;
    end

    assign uInstruction = uInstructionStore[uPC];

endmodule
